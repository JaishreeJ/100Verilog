module demux1_4_tb;
wire [3:0] Y;
reg [1:0] A;
reg din;
demux1_4 demux (Y, A, din);
initial begin
    din = 1;
    A = 2'b00;
#1  A = 2'b01;
#1  A = 2'b10;
#1  A = 2'b11;
end
initial begin
    $monitor("%t| Din = %d| A[1] = %d| A[0] = %d| Y[0] = %d| Y[1] = %d| Y[2] = %d| Y[3] = %d",
              $time, din, A[1], A[0], Y[0], Y[1], Y[2], Y[3]);
  $dumpfile("dump.vcd");
  $dumpvars(1);
end
endmodule
